`include "hello_world/hello_world.v"
module module_call;

endmodule
