module dflipflop (clk,din, dout);

input wire clk, din;

output dout;

always @(posclk)
//define d flipflop

endmodule