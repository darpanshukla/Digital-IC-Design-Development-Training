// ref: https://github.com/yasnakateb/WMController
`include "Microcontroller.v"
module Microcontroller_tb();
    reg clock;
    reg input1;
    reg input2;
    reg input3;
    reg input4;
    reg input5;
    reg input6;
    reg sig_Lid_Closed;
    reg sig_Coin;
    reg sig_Cancel;
    reg sig_Time_Out;
    reg sig_Out_Of_Balance;
    reg sig_Motor_Failure;
    wire [2:0] state;

Microcontroller uut(
    .clock(clock),
    .input1(input1),
    .input2(input2),
    .input3(input3),
    .input4(input4),
    .input5(input5),
    .input6(input6),
    .sig_Lid_Closed(sig_Lid_Closed),
    .sig_Coin(sig_Coin),
    .sig_Cancel(sig_Cancel),
    .sig_Time_Out(sig_Time_Out),
    .sig_Out_Of_Balance(sig_Out_Of_Balance),
    .sig_Motor_Failure(sig_Motor_Failure),
    .state(state)
    );

    always #1 clock = ~ clock;

    initial begin 
    $dumpfile("Microcontroller_tb.vcd");
    $dumpvars(0,Microcontroller_tb);

        clock = 0;
        sig_Coin = 1;
        sig_Lid_Closed = 1;
        input1 = 0;
        input2 = 1;
        input3 = 0;
        input4 = 0;
        input5 = 0;
        input6 = 0;

        #100
        input2 = 0;
        input6 = 1;
    end

    initial #1000 $finish;

endmodule
