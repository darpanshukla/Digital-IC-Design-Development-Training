module top_level_baud_rate_generator_tb;

// Instantiate the Testbench for Baud Rate Generator module
testbench_baud_rate_generator tb();

endmodule
